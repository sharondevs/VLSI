module port_assignment_stage1(output reg port_num,input [31:0]flit);
	always@(*)begin
	case(flit[6:4])
	3'b000 : port_num = 0;
	3'b001 : port_num = 1;
	3'b010 : port_num = 0;
	3'b011 : port_num = 1;
	endcase 
end
endmodule

module exchanger_stage1(output reg[31:0] flit_0_out,flit_1_out, input prio_flit_num, input [31:0]flit_0,flit_1);
	reg [31:0] prio_flit;
	reg stage = 0;
	wire port_num;
	port_assignment_stage1 assign_block1(.port_num(port_num), .flit(prio_flit));
	always@(*)begin
	if(prio_flit_num == 0)begin
	prio_flit = flit_0;
		if(port_num == 0) begin
		flit_0_out = prio_flit;
		flit_1_out = flit_1;
		end
		else begin
		flit_1_out = prio_flit;
		flit_0_out = flit_1;
		end
	end else begin
	prio_flit = flit_1;
		if(port_num == 0) begin
		flit_0_out = prio_flit;
		flit_1_out = flit_0;
		end else begin
		flit_1_out = prio_flit;
		flit_0_out = flit_0;
		end
	end
end
endmodule


module permuter_stage1(output [31:0] per_out_0,per_out_1 ,input [31:0] per_in_0,per_in_1 );
	wire sel_flit_num;
	arbiter arb(.winner(sel_flit_num), .arb_in_0(per_in_0), .arb_in_1(per_in_1));
	exchanger_stage1 exchange(.prio_flit_num(sel_flit_num),.flit_0(per_in_0), .flit_1(per_in_1), .flit_0_out(per_out_0), .flit_1_out(per_out_1));
endmodule 

module port_assignment_stage2(output reg port_num,input [31:0]flit);
	always@(*)begin
	case(flit[6:4])
	3'b000 : port_num = 0;
	3'b001 : port_num = 0;
	3'b010 : port_num = 1;
	3'b011 : port_num = 1;
	endcase 
end
endmodule

module exchanger_stage2(output reg [31:0] flit_0_out,flit_1_out, input prio_flit_num, input [31:0]flit_0,flit_1);
	reg [31:0] prio_flit;
	reg stage = 0;
	wire port_num;
	port_assignment_stage2 assign_block2(.port_num(port_num), .flit(prio_flit));
	always@(*)begin
	if(prio_flit_num == 0)begin
	prio_flit = flit_0;
		if(port_num == 0) begin
		flit_0_out = prio_flit;
		flit_1_out = flit_1;
		end
		else begin
		flit_1_out = prio_flit;
		flit_0_out = flit_1;
		end
	end else begin
	prio_flit = flit_1;
		if(port_num == 0) begin
		flit_0_out = prio_flit;
		flit_1_out = flit_0;
		end else begin
		flit_1_out = prio_flit;
		flit_0_out = flit_0;
		end
	end
end
endmodule

module permuter_stage2(output [31:0] per_out_0,per_out_1 ,input [31:0] per_in_0,per_in_1 );
	wire sel_flit_num;
	arbiter arb(.winner(sel_flit_num), .arb_in_0(per_in_0), .arb_in_1(per_in_1));
	exchanger_stage2 exchange(.prio_flit_num(sel_flit_num),.flit_0(per_in_0), .flit_1(per_in_1), .flit_0_out(per_out_0), .flit_1_out(per_out_1));
endmodule 

/*
The block instantiations in the permuter engine corresponds to the different arbiters in the permutation block
Block1 - The upper block in stage 1 (N,E inputs)
Block2 - The lower block in stage 1 (S,W inputs)
Block3 - The upper block in stage 2
Block4  - The lower block in stage 2
*/
module permutation_engine(output [31:0] PNout,PEout, PSout,PWout, input [31:0] PNin,PEin,PSin,PWin); 
	wire [31:0]inter_con1,inter_con2, inter_con3,inter_con4;
	// Stage 1 -
	permuter_stage1 block1(.per_out_0(inter_con1),.per_out_1(inter_con2) ,.per_in_0(PNin),.per_in_1(PEin));
	permuter_stage1 block2(.per_out_0(inter_con3),.per_out_1(inter_con4) ,.per_in_0(PSin),.per_in_1(PWin));
	// Stage 2 -
	permuter_stage2 block3(.per_out_0(PNout),.per_out_1(PSout) ,.per_in_0(inter_con1),.per_in_1(inter_con3));
	permuter_stage2 block4(.per_out_0(PEout),.per_out_1(PWout) ,.per_in_0(inter_con2),.per_in_1(inter_con4));

endmodule
